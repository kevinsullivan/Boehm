(** ** STAGE MODULE *)
(**
Kevin Sullivan, Chong Tang, Ke Dou, with Donna Rhodes, 
Barry Boehm, and Adam Ross 

March, 2015
*)

(** 
This module defines the [Stage], which represents the stages (or processes) 
that the system needs to be involved in.
*)
Module Stage.
  Inductive Stage := aStage.
End Stage.
